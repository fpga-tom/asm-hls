/*
* This is full adder
*/

module full_adder
(
	input x,
	input y,
	output z
);

assign z = x + y;

endmodule
